LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Calc IS
    PORT( 
        A_bin       : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        B_bin       : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
        Add_Or_Mul  : IN  STD_LOGIC;
        Sum_Or_Sub  : IN  STD_LOGIC;
        Result      : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
    );
END ENTITY Calc;

ARCHITECTURE behaviour OF Calc IS

	 SIGNAL A_Sum_Sub      : STD_LOGIC_VECTOR(4 DOWNTO 0);
	 SIGNAL B_Sum_Sub      : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL Add_Sub_Result : STD_LOGIC_VECTOR(4 DOWNTO 0);
    SIGNAL Add_Sub_Ext    : STD_LOGIC_VECTOR(6 DOWNTO 0);
    SIGNAL Mul_Result     : STD_LOGIC_VECTOR(6 DOWNTO 0);
    SIGNAL Cout_Sign      : STD_LOGIC;

BEGIN

	A_Sum_Sub <= "0" & A_bin;
	B_Sum_Sub <= "0" & B_bin;

   Add_Sub: ENTITY work.N_Adder
        GENERIC MAP (
            N => 5
        )
        PORT MAP(
            ina  => A_Sum_Sub,
            inb  => B_Sum_Sub,
            sign => Sum_Or_Sub,
            sum  => Add_Sub_Result,
            Cout => Cout_Sign
        );

    Mul: ENTITY work.Mult4x7
        PORT MAP(
            a    => A_Bin,
            b    => B_Bin,
            prod => Mul_Result
        );

    Add_Sub_Ext <= "00" & Add_Sub_Result WHEN Cout_Sign = '1' ELSE "11" & Add_Sub_Result;

    Result <= Add_Sub_Ext WHEN Add_Or_Mul = '1' ELSE Mul_Result;

END behaviour;
